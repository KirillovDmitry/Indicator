`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// ������ ����������� ��������� ����� �� �������������� ����������.
// ��������� ����������� ������������������ �������� �����, ������� ������������ �� ����������.
// ����������� ��� �������� �������: ���� �������������� ���������� ��������� ����������, ������ 
// �������������� ������������ ��������� �������� �������� ������.
//
//////////////////////////////////////////////////////////////////////////////////

module main(

    input  tg, // ������� �������� ������� � ������ (�� ���������� ����� f = 25���)
    
	output S1, // ������ ������ �������� ������� ����������
    output S2, // 
    output S3, // 
    output S4, // ������ ������ �������� ������� ����������
	
    output DA, // ��������� �������� ���������� // 7-segment encoding
    output DB, // ��������� �������� ���������� //      0
    output DC, // ��������� �������� ���������� //     ---
    output DD, // ��������� �������� ���������� //  5 |   | 1
    output DE, // ��������� �������� ���������� //     --- <--6
    output DF, // ��������� �������� ���������� //  4 |   | 2
    output DG  // ��������� �������� ���������� //     ---
    											//      3
);

	//-----------------------------------------------------------	
	// �������� ������� �������
	always @(posedge tg)
			REG <= REG + 1'b1; 
	
	parameter par = 15;
	reg [25:0] REG = 0;
	reg clc = 0;
	always @(posedge REG[par])
		clc = ~clc;
		
	//-----------------------------------------------------------	
	// ������������ �������� ������
	reg [13:0] D_ = 0;		
	always @(negedge REG[par+3])
		if (D_ < 9999)
			D_ <= D_ + 1'b1;
		else 
			D_ = 0;
		
	//-----------------------------------------------------------	
	// �������� ������ �������-����������� �������������� ������
	// � ������ �� �� ������������ ���������
	wire [13:0] D;
	wire [17:0] Q;			
	assign D = D_;
	BinToInd uut3(.D(D), .tg(clc), .S1(S1), .S2(S2), .S3(S3), .S4(S4), .DA(DA), .DB(DB), .DC(DC), .DD(DD),
    .DE(DE), .DF(DF), .DG(DG) );

endmodule
