`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// ������ ������������� �������-����������� ��������������
//
//////////////////////////////////////////////////////////////////////////////////

module EP(
    input  [3:0] X,
    output [3:0] Y
);

assign Y = (X<=4)? X : X + 4'd3;

endmodule
