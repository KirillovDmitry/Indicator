`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// ������ �������������� ��������� ���� � �������-���������� (���8421) ���.
// �������������� �������������� ������������� �������, ��������� � 
// ����� �., ���� �. ����������������� ������������: ���������� ����������� �� ��� 323 ���� 19.6
// ����� ����� ��� �������������� ������������ ���������������� ��������� ���������.
//
//////////////////////////////////////////////////////////////////////////////////

module BinToDec8421(
    input  [13:0] D, // ������� �������, ���������� �������� ���
    output [17:0] Q	 // �������� �������, ���������� ���8421
);
	// �������� ���������� �������������� ����������
	wire [3:0]  Q1;
	wire [3:0]  Q2;
	wire [3:0]  Q3;
	wire [7:0]  Q4;
	wire [7:0]  Q5;
	wire [7:0]  Q6;
	wire [11:0] Q7;
	wire [11:0] Q8;
	wire [11:0] Q9;
	wire [14:0] Q10;

	// �������������� �������������� ����� ���������������-�������������
	// ����������� ������� ������������� �������������� EP
	EP uut1 (
			.X({1'b0, D[13:11]}), 
			.Y(Q1[3:0])
		);
	
	//-------------------------	

	EP uut2 (
			.X({Q1[2:0], D[10]}), 
			.Y(Q2[3:0])
		);
		
	//-------------------------		

	EP uut3 (
			.X({Q2[2:0], D[9]}), 
			.Y(Q3[3:0])
		);	
		
	//-------------------------	

	EP uut4 (
			.X({1'b0, Q1[3], Q2[3], Q3[3]}), 
			.Y(Q4[7:4])
		);	

	EP uut5 (
			.X({Q3[2:0], D[8]}), 
			.Y(Q4[3:0])
		);	
		
	//-------------------------	

	EP uut6 (
			.X({Q4[6:3]}), 
			.Y(Q5[7:4])
		);	

	EP uut7 (
			.X({Q4[2:0], D[7]}), 
			.Y(Q5[3:0])
		);	
		
	//-------------------------	

	EP uut8 (
			.X(Q5[6:3]), 
			.Y(Q6[7:4])
		);	

	EP uut9 (
			.X({Q5[2:0], D[6]}), 
			.Y(Q6[3:0])
		);		
		
	//-------------------------	

	EP uut10 (
			.X({1'b0, Q4[7], Q5[7], Q6[7]}), 
			.Y(Q7[11:8])
		);	

	EP uut11 (
			.X(Q6[6:3]), 
			.Y(Q7[7:4])
		);

	EP uut12 (
			.X({Q6[2:0], D[5]}), 
			.Y(Q7[3:0])
		);		
		
	//-------------------------	

	EP uut13 (
			.X(Q7[10:7]), 
			.Y(Q8[11:8])
		);	

	EP uut14 (
			.X(Q7[6:3]), 
			.Y(Q8[7:4])
		);

	EP uut15 (
			.X({Q7[2:0], D[4]}), 
			.Y(Q8[3:0])
		);		
		
	//-------------------------	

	EP uut16 (
			.X(Q8[10:7]), 
			.Y(Q9[11:8])
		);	

	EP uut17 (
			.X(Q8[6:3]),
			.Y(Q9[7:4])
		);

	EP uut18 (
			.X({Q8[2:0], D[3]}), 
			.Y(Q9[3:0])
		);	
		
	//-------------------------	

	EP uut19 (
			.X({1'b0, Q7[11], Q8[11], Q9[11]}), 
			.Y({Q[17], Q10[14:12]})
		);	
		
	EP uut20 (
			.X(Q9[10:7]), 
			.Y(Q10[11:8])
		);	

	EP uut21 (
			.X(Q9[6:3]), 
			.Y(Q10[7:4])
		);

	EP uut22 (
			.X({Q9[2:0], D[2]}), 
			.Y(Q10[3:0])
		);		
		
	//-------------------------	

	EP uut23 (
			.X(Q10[14:11]), 
			.Y(Q[16:13])
		);	
		
	EP uut24 (
			.X(Q10[10:7]), 
			.Y(Q[12:9])
		);	

	EP uut25 (
			.X(Q10[6:3]), 
			.Y(Q[8:5])
		);

	EP uut26 (
			.X({Q10[2:0], D[1]}), 
			.Y(Q[4:1])
		);		
		
	//-------------------------	

	// ������� Q �������� �������� ��������� ��������������
	assign Q[0] = D[0];

endmodule
