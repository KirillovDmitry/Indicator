`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// ������ ������ ��������� ��������� �������� �� ��������� ���������� �����
//
//////////////////////////////////////////////////////////////////////////////////

module BinToInd(
    input  [13:0] D,		// ������� ������� �������� ������ ��� ����������� �� ����������
    input  tg, 			    // ������� ���������� ����������
    output S1,				// ������ ������ ������� �������� ����������
    output S2,				// ������ ������ ������� �������� ����������
    output S3,				// ������ ������ �������� �������� ����������
    output S4,				// ������ ������ ���������� �������� ����������
    output DA,				// ��������� �������� ���������� // 7-segment encoding
    output DB,				// ��������� �������� ���������� //      0
    output DC,				// ��������� �������� ���������� //     ---
    output DD,				// ��������� �������� ���������� //  5 |   | 1
    output DE,				// ��������� �������� ���������� //     --- <--6
    output DF,				// ��������� �������� ���������� //  4 |   | 2
    output DG				// ��������� �������� ���������� //     ---
);														     //      3

	//-----------------------------------------------------------
	// ������� ������ �������� ������ ����������� � ������� ���������� ��� ���8421
	wire [17:0] Q;
	BinToDec8421 uut ( .D(D), .Q(Q) );
	
	// ���������� NumInd �������� ���� ������� ������� ���������� ��� �����������,
	// ��������� �������� �� ���������� �, �������������, ������
	reg [1:0] NumInd = 0;
	always @(posedge tg)
		NumInd <= NumInd + 1'b1;
		
	// S_SEG ��������� ������ ������ �������� ��������, � Dec8421 ������������
	// ������ �������� ��� ��� ������ �� ������� ������� ����������
	reg [3:0] S_SEG = 0;
	reg [3:0] Dec8421 = 0;
	always @(negedge tg)
		case (NumInd)
			 2'b00 : begin S_SEG = 4'b1000; Dec8421 = Q[3:0];   end
			 2'b01 : begin S_SEG = 4'b0100; Dec8421 = Q[7:4];   end
			 2'b10 : begin S_SEG = 4'b0010; Dec8421 = Q[11:8];  end
			 2'b11 : begin S_SEG = 4'b0001; Dec8421 = Q[16:12]; end
		endcase
	
	// �������� ��������, ����������� ��� ��� ������ �� ������� ������� ��������
	// ������������� � ���������� ��� ��������� �����������
	wire [6:0] IND;		
	DecToInd uut (.Dec(Dec8421),.Ind(IND));	
	
	//-----------------------------------------------------------	
	// �� �������� �������� ������� ������� ������ �������� �������� � ������� ���������
	// ��������� �����������
	assign S1 = ~S_SEG[0];
	assign S2 = ~S_SEG[1];
	assign S3 = ~S_SEG[2];
	assign S4 = ~S_SEG[3];

	assign DA = IND[0];
	assign DB = IND[1];
	assign DC = IND[2];
	assign DD = IND[3];
	assign DE = IND[4];
	assign DF = IND[5];
	assign DG = IND[6];

endmodule
